module aish_inverter(output Y, input A);
    not (Y, A);
endmodule